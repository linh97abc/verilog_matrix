module add__ (
    input clk,
    input reset,
    input clk_en,
    input [31:0] a,
    input [31:0] b,
    output [31:0] q,
    input start,
    output wire done
);
    
endmodule