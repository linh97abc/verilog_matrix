module custom_instruct (
    input [31:0] dataa,
    input [31:0] datab,
    input [31:0] result,
    input clk,
    input clk_en,
    input start,
    input reset,
    output done,
    input [7:0] n
);
    
endmodule